module part2_64_tb();

		logic [63:0] x, y;
		logic [63:0] result;

		logic zero, underflow, overflow, nan;

		part2 #(.E(11), .M(52)) DUT (
			.X(x),
			.Y(y),
			.result(result),
			.zero(zero),
			.underflow(underflow),
			.overflow(overflow),
			.nan(nan)
		);


		initial begin
			// Testing normal operation
			// 224.5*-254.78
			x = 64'b0100000001101100000100000000000000000000000000000000000000000000;
			y = 64'b1100000001101111110110001111010111000010100011110101110000101001;
			#10;
			if (result != 64'b1100000011101011111011011100001110000101000111101011100001010001) begin
				$display("Error! 224.5*-254.78");
				$stop();
			end

			// -433.24 * -4.5
			x = 64'b1100000001111011000100111101011100001010001111010111000010100100;
			y = 64'b1100000000010010000000000000000000000000000000000000000000000000;
			#10;
			if (result != 'b0100000010011110011101100101000111101011100001010001111010111000) begin
				$display("Error! -433.24 * -4.5");
				$stop();
			end



			//Special Case
			//Zero
			// +zero * #!=inf	->E=0,M=0,zero=1
			x = 64'b0;
			y = 64'b0100000000010010000000000000000000000000000000000000000000000000;
			#10;
			if (result != 64'b0 || zero == 1'b0) begin
				$display("Error! zero1");
				$stop();
			end


			// #!=inf * -zero	->E=0,M=0,zero=1
			x = 64'b0000000000000000000000000000000000000000000000000000000000000000;
			y = 64'b1100000000010010000000000000000000000000000000000000000000000000;
			#10;
			if (result != 64'b1000000000000000000000000000000000000000000000000000000000000000 || zero == 1'b0) begin
				$display("Error! zero1");
				$stop();
			end

			//NaN
			// +zero * #=inf	->S=0, E=EB,M=0,NaN=1
			x = 64'b0 ;
			y = 64'b0111111111111010101001001100110100000101001010010010101010010010;
			#10;
			if (result != 64'b0111111111110000000000000000000000000000000000000000000000000000||nan==1'b0) begin
				$display("Error! NaN1");
				$stop();
			end

			// #=-inf * zero	->S=1, E=EB,M=0,Nah=1
			x = 64'b1111111111110101101011010010101010010010010011100000000000000000;
			y = 64'b0100000100011000000100100111101001010001010000100100101001010010;
			#10;
			if (result != 64'b1111111111110000000000000000000000000000000000000000000000000000||nan==1'b0) begin
				$display("Error! NaN2");
				$stop();
			end

			//Underflow
			//s=0, E <0	->E=0,M!=0,underflow=1
			x = 64'b0000010000010100110000000000000000000000110000000000000000000000;
			y = 64'b0001000100011001100000000000000000000000000100100111010100101001;
			#10;
			if (result != 64'b0000000000000000000000000000000000000000000000000000000000000001 || underflow == 0) begin
				$display("Error! Underflow1");
				$stop();
			end

			//s=1, E <0	->E=0,M!=0,underflow=1
			x = 64'b0000010000010100110000000000000000000000110000000001100000000100;
			y = 64'b0000000100101001100000000000000000000001100000000000000100000000;
			#10;
			if (result != 64'b0000000000000000000000000000000000000000000000000000000000000001 || underflow == 0) begin
				$display("Error! Underflow2");
				$stop();
			end

			//overflow
			// E >= 2**(E)-1, 2**(E)-1, M=0, overflow=1
			x = 64'b1111110111111011100000000001010100101001010101010001001001010101;
			y = 64'b1111101111110000000001000010000101010101001010011010100100010101;
			#10;
			if (result != 64'b0111111111110000000000000000000000000000000000000000000000000000 || overflow == 1'b0) begin
				$display("Error! Overflow2");
				$stop();
			end



			$display("The test passed");
			$stop();
		end
endmodule
